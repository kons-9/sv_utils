`ifndef COLOR_SVH
`define COLOR_SVH

`include "color_impl.svh"

`define BLACK_COLOR `BLACK_COLOR_IMPL
`define RED_COLOR `RED_COLOR_IMPL
`define GREEN_COLOR `GREEN_COLOR_IMPL 
`define YELLOW_COLOR `YELLOW_COLOR_IMPL
`define BLUE_COLOR `BLUE_COLOR_IMPL
`define MAGENTA_COLOR `MAGENTA_COLOR_IMPL
`define CYAN_COLOR `CYAN_COLOR_IMPL
`define WHITE_COLOR `WHITE_COLOR_IMPL
`define GRAY_COLOR `GRAY_COLOR_IMPL
`define RESET_COLOR `RESET_COLOR_IMPL

`endif
