`ifndef SV_TEST_IMPL_SVH
`define SV_TEST_IMPL_SVH

`define TEST_SECTION_START_IMPL(section_name)
`define ENABLE_FATAL_IMPL()
`define DISABLE_FATAL_IMPL()
`define TEST_START_IMPL(test_log_path)
`define TEST_EXPECTED_IMPL(expected, actual, message, file, line)
`define TEST_UNEXPECTED_IMPL(unexpected, actual, message, file, line)
`define TEST_RESULT_IMPL()

`endif
