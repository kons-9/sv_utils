`define DISABLE_FATAL_EXIT_IMPL
