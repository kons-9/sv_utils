`ifndef LOG_IMPL_SVH
`define LOG_IMPL_SVH

`define LOG_IMPL(level, tag, msg, file, line)
`define LOG_VERBOSE_IMPL(tag, msg)
`define LOG_DEBUG_IMPL(tag, msg)
`define LOG_INFO_IMPL(tag, msg)
`define LOG_WARN_IMPL(tag, msg)
`define LOG_ERROR_IMPL(tag, msg)
`define LOG_FATAL_IMPL(tag, msg)

`endif
