`ifndef EXIT_SVH
`define EXIT_SVH

`include "exit_impl.svh"

`define DISABLE_FATAL_EXIT `DISABLE_FATAL_EXIT_IMPL

`endif
